`timescale 1ns / 1ps

/*******************************************************************
*
* Module: InstMem.v
* Project: Milestone 2
* Author: Mohamed Abbas mohamed_abbas02@aucegypt 
          Omar Bahgat omar_bahgat@aucegypt.edu
* Description: Instruction Memory
*
* Change history: 
**********************************************************************/

module InstMem (
    input [5:0] addr, 
    output [31:0] data_out
); 
    
   reg [31:0] mem [0:63];
   initial begin
   
        // R-format Instructions
        
        mem[0]=32'b000000000000_00000_010_00001_0000011 ; //lw x1, 0(x0) 10
        mem[1]=32'b000000000100_00000_010_00010_0000011 ; //lw x2, 4(x0) 5
        mem[2]=32'b0000000_00010_00001_000_00011_0110011 ; //add x3, x1, x2 15
        mem[3]=32'b0100000_00010_00001_000_01000_0110011 ; //sub x8, x1, x2 5
        mem[4]=32'b0000_0000_0010_0000_1100_0010_1011_0011;   // xor x5, x1, x2 15
        mem[5] =32'b0000_0000_0010_0000_1110_0011_0011_0011;   // or x6, x1, x2
        mem[6] = 32'b001000001111001110110011;   // and x7, x1, x2
        mem[7] = 32'b0010_0000_1001_0100_0011_0011;   // sll x8, x1, x2
        mem[8] = 32'b001000001101010010110011;   // srl x9, x1, x2
        mem[9] = 32'b01000000001000001101010100110011;   // sra x10, x1, x2

//        mem[10] = 8'h0020a5b3;  // slt x11, x1, x2
//        mem[11] = 8'h0020b633;  // sltu x12,x1, x2

          // I-format Instructions

//        mem[2] = 32'b010000001000010100010011;  // addi x10, x1, 4
//        mem[3] = 32'b010000001100010100010011;  // xori x10, x1, 4
//        mem[4] = 32'b010000001110010100010011;// ori x10, x1, 4
//        mem[5] = 32'b010000001111010100010011;// andi x10, x1, 4
//        mem[6] = 32'b010000001001010100010011;// slli x10, x1, 4
//        mem[7] = 32'b010000001101010100010011;// srli x10, x1, 4
//        mem[8] = 32'b01000000010000001101010100010011;// srai x10, x1, 4

//        mem[9] = 32'b010000001010010100010011;// slti x10, x1, 4
//        mem[10] = 32'b010000001011010100010011;// sltiu x10, x1, 4

        // Load Instructions

//        mem[2] = 32'b000110000011;      // lb x3, 0(x0)
//        mem[3] = 32'b0001000110000011;  // lh x3, 0(x0)
//        mem[4] = 32'b0010000110000011;  // lw x3, 0(x0)
//        mem[5] = 32'b0100000110000011;  // lbu x3, 0(x0)
//        mem[6] = 32'b0101000110000011;  // lhu x3, 0(x0)


        // Store Instructions 
        
//        mem[2] = 32'b000100000000000000100011;  // sb x1, 0(x0)
//        mem[3] = 32'b000100000001000000100011;  // sh x1, 0(x0)
//        mem[4] = 32'b000100000010000000100011;  // sw x1, 0(x0)
        
//        // Branch Instructions
        
//        mem[2] = 32'b1000010001100011;          // beq x0, x0, 8
        
//        mem[3] = 32'b000100000000000110010011;  // add x3, x0, 1
//        mem[4] = 32'b001000000000000110010011;  // add x3, x0, 2
        
//        mem[5] = 32'b0001010001100011;          // bne x0, x0, 8
        
//        mem[6] = 32'b000100000000000110010011;
//        mem[7] = 32'b001000000000000110010011;
        
//        mem[8] = 32'b0100010001100011;          // blt x0, x0, 8
        
//        mem[9] = 32'b000100000000000110010011;
//        mem[10] = 32'b001000000000000110010011;
        
//        mem[11] = 32'b0101010001100011;         // bge x0, x0, 8
        
//        mem[12] = 32'b000100000000000110010011;
//        mem[13] = 32'b001000000000000110010011;
        
//        mem[14] = 32'b0110010001100011;         // bltu x0, x0, 8
        
//        mem[15] = 32'b000100000000000110010011;
//        mem[16] = 32'b001000000000000110010011;
        
//        mem[17] = 32'b0111010001100011;         // bgeu x0, x0, 8

//        mem[18] = 32'b000100000000000110010011;
//        mem[19] = 32'b001000000000000110010011;
        
    end
    assign data_out = mem[addr]; 
endmodule