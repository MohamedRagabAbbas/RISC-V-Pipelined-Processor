`timescale 1ns / 1ps

/*******************************************************************
*
* Module: InstMem.v
* Project: Milestone 2
* Author: Mohamed Abbas mohamed_abbas02@aucegypt 
          Omar Bahgat omar_bahgat@aucegypt.edu
* Description: Instruction Memory
*
* Change history: 
**********************************************************************/

module InstMem (
    input [5:0] addr, 
    output [31:0] data_out
); 
    
   reg [31:0] mem [0:63];
   initial begin
   
        mem[0] = 8'h00002083;   // lw x1, 0(x0)
        mem[1] = 8'h00402103;   // lw x2, 4(x0)
        mem[2] = 8'h002081b3;   // add x3, x1, x2
        mem[3] = 8'h40208233;   // sub x4, x1, x2
        mem[4] = 8'h0020c2b3;   // xor x5, x1, x2
        mem[5] = 8'h0020e333;   // or x6, x1, x2
        mem[6] = 8'h0020f3b3;   // and x7, x1, x2
        mem[7] = 8'h00209433;   // sll x8, x1, x2
        mem[8] = 8'h0020d4b3;   // srl x9, x1, x2
        mem[9] = 8'h4020d533;   // sra x10, x1, x2
        mem[10] = 8'h0020a5b3;  // slt x11, x1, x2
        mem[11] = 8'h0020b633;  // sltu x12,x1, x2

//        mem[0]=32'b000000000000_00000_010_00001_0000011 ; //lw x1, 0(x0) 17
//        mem[1]=32'b000000000100_00000_010_00010_0000011 ; //lw x2, 4(x0) 9 
//        mem[2]=32'b000000001000_00000_010_00011_0000011 ; //lw x3, 8(x0) 25 
//        mem[3]=32'b0000000_00010_00001_110_00100_0110011 ; //or x4, x1, x2 25
//        mem[4]=32'b0_000000_00011_00100_000_0100_0_1100011; //beq x4, x3, 0
//        mem[5]=32'b0000000_00010_00001_000_00011_0110011 ; //add x3, x1, x2 
//        mem[6]=32'b0000000_00010_00011_000_00101_0110011 ; //add x5, x3, x2 34
//        mem[7]=32'b0000000_00101_00000_010_01100_0100011; //sw x5, 12(x0) x
//        mem[8]=32'b000000001100_00000_010_00110_0000011 ; //lw x6, 12(x0)  34
//        mem[9]=32'b0000000_00001_00110_111_00111_0110011 ; //and x7, x6, x1 addr
//        mem[10]=32'b0100000_00010_00001_000_01000_0110011 ; //sub x8, x1, x2 8
//        mem[11]=32'b0000000_00010_00001_000_00000_0110011 ; //add x0, x1, x2 x
//        mem[12]=32'b0000000_00001_00000_000_01001_0110011 ; //add x9, x0,x1 addr 17
    end
    assign data_out = mem[addr]; 
endmodule